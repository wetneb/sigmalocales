
(** Formalization of Theorem 3.3 in 
  
   Thierry Coquand, Giovanni Sambin, Jan Smith, Silvio Valentini

   Inductively generated formal topologies

   #<a href="http://doai.io/10.1016/S0168-0072(03)00052-6">http://doai.io/10.1016/S0168-0072(03)00052-6</a>#
 
   Adapted to distributive lattices. See
   the [FreeFrame] module for more insightful comments
   (this is the same proof, just for finite formal joins
    instead of countable ones). I have some ideas about
   how to refactor the two in the same proof: define the free 
   kappa-frame generated by a meet semilattice with axioms,
   where kappa is the appropriate constructive cardinal-like 
   object…

 *)

Require Import MathClasses.interfaces.canonical_names.
Require Import BijNat.
Require Import Frame.
Require Import MeetSemiLattice.
Require Import PreorderEquiv.
Require Import DistrLattice.
Require Import Coq.Classes.RelationClasses.
Require Import Coq.Lists.List.
Require Import Coq.Lists.SetoidList.

Section Definition_Inductive_Locale.

  (** * Definition of the free distributive lattice *)
  
  (** Generators. *)
  Variable T : Type.
  Variable Tle : Le T.
  Variable Tmsl : @MeetSemiLattice T Tle.
  Existing Instance Tmsl.
  Existing Instance Feq_equiv.
  Existing Instance Feq_equivalence.
 
  (** For each generator, an index set for its coverings. *)
  Variable Idx : forall t:T, Set.
  (** For each generator and index of covering, an covering. *)
  Variable CovAx : forall t:T, forall i:Idx t, list T.
  
  (** ** Preliminaries on finite sets with lists *)
  
  Notation "( a ⊓)" := (fun el => a ⊓ el).
  
  Definition down (a : T) (U : list T) : list T :=
    map (a ⊓) U.

  Infix "↓" := down (at level 50).

  Infix "↪" := (inclA Feq) (at level 75).
  Instance in_contains : Contains T (list T) := (InA Feq).

  Lemma inclA_app_l : forall u v, u ↪ u ++ v.
  Proof.
    unfold inclA ; intros.
    rewrite InA_app_iff.
    left. assumption.
  Qed.

  Lemma inclA_app_r : forall u v, v ↪ u ++ v.
  Proof.
    unfold inclA ; intros.
    rewrite InA_app_iff.
    right. assumption.
  Qed.

  Lemma map_in : forall f x U, (Proper ((=) ==> (=)) f) -> x ∈ U -> f x ∈ map f U.
  Proof.
    intros. unfold map.
    induction H0.
    apply InA_cons_hd.
    apply H. assumption.
    apply InA_cons_tl.
    assumption.
  Qed.

  Lemma in_map : forall f x U, x ∈ map f U -> exists y, y ∈ U /\ x = f y.
  Proof.
    intros.
    induction U.
    - inversion H.
    - set (V := map f (a :: U)) in *. assert( V ≡ map f (a :: U)) by reflexivity.
      destruct H.
      + inversion H0.
        exists a. split.
        apply InA_cons_hd. reflexivity.
        rewrite <- H2. assumption.
      + simpl in H0.
        inversion H0. subst.
        apply IHU in H.
        destruct H as [y [G K]].
        exists y. split.
        apply InA_cons_tl.
        assumption. assumption.
  Qed.

  Instance FeqT_equivalence : Equivalence (Feq : T -> T -> Prop).
  Proof.
    apply Feq_equivalence.
    apply (@msl_preorder T le Tmsl).
  Qed.

  Instance InA_Feq_compat : Proper (Feq ==> equivlistA Feq ==> iff) (InA (Feq : Equiv T)) := (InA_compat FeqT_equivalence).

  Definition equiv_listT : list T -> list T -> Prop := equivlistA Feq.
  Add Setoid (list T) equiv_listT (equivlist_equiv FeqT_equivalence) as equiv_listT_setoid.
  Infix "==" := equiv_listT (at level 75).

  (** ** Inductive cover relation
   Here, we need an additional axiom to equate [[]] and
   [[⊥]].
   *)
  
  Inductive covrel (a : T) : (list T) -> Prop :=
  | cr_bot : forall U, a = ⊥ -> covrel a U
  | cr_refl : forall U, a ∈ U -> covrel a U
  | cr_inf : forall U b, forall i:Idx b, a ≤ b -> (forall x, x ∈ (CovAx b i) -> covrel (a ⊓ x) U) -> covrel a U
  | cr_left : forall U b, a ≤ b -> covrel b U -> covrel a U.
  Infix "◁" := (covrel) (at level 60).

  Lemma covrel_Teq : forall x: T, forall U, (x ◁ U) -> forall y :T,  x = y -> y ◁ U.
  Proof.
    intros.
    destruct H0.
    apply cr_left with (b := x) ; assumption.
  Qed.
    
  Lemma covrel_proper : Proper ((=) ==> eq ==> iff) covrel.
  Proof.
    unfold Proper, respectful.
    intros.
    split ; intro.
    
    rewrite <- H0.
    apply (covrel_Teq x x0 H1 y H).

    rewrite H0.
    apply (covrel_Teq y y0 H1 x).
    symmetry. apply H.
  Qed.
  Add Parametric Morphism : covrel with signature ((=) ==> eq ==> iff) as covrel_morphism.
  Proof.
    intros. apply covrel_proper. apply H. reflexivity.
  Qed.

  (** ** Preorder and equivalence between coverings *)

  Definition Covrel (U V : list T) :=
    forall x, x ∈ U -> x ◁ V.
  Instance Covrel_le : Le (list T) := Covrel.
  Ltac unfold_Covrel := unfold le, Covrel_le, Covrel.
  Ltac unfold_Covrel_in a := unfold le, Covrel_le, Covrel in a.

  
  Lemma cr_trans : forall (a : T) (U W : list T), a ◁ U -> U ≤ W -> a ◁ W.
  Proof.
    intros a U W CR.
    generalize W ; clear W.
    induction CR ; intros.
    - (* cr_bot *)
      destruct W.
      apply cr_bot ; assumption.
      apply cr_left with (b := t).
      rewrite H. apply bot_le.
      apply cr_refl. apply InA_cons_hd. reflexivity.
    - (* cr_refl *)
      unfold_Covrel_in H0.
      apply H0. assumption.
    - (* cr_inf *)
      apply (cr_inf a W b i H).
      intros. apply H1 ; assumption.
    - (* cr_left *)
      apply cr_left with (b := b).
      assumption.
      apply IHCR ; apply H0.
  Qed.

  Lemma Covrel_refl : Reflexive Covrel.
  Proof.
    unfold Reflexive.
    intros.
    unfold Covrel.
    intros. apply cr_refl.
    assumption.
  Qed.
    
  Lemma Covrel_trans : Transitive Covrel.
  Proof.
    unfold Transitive, Covrel.
    intros.
    apply cr_trans with (U := y).
    apply H. assumption.
    assumption.
  Qed.

  Definition PO_for_FDistrLattice : @Preorder (list T) Covrel :=
    MkPreorder
      (list T)
      Covrel
      Covrel_refl
      Covrel_trans.
  Existing Instance PO_for_FDistrLattice.
  
  Add Morphism covrel : covrel_morphism2.
  Proof.
    intros x y Heq U W H.
    destruct H as [Hl Hr].
    split ; intro.
    apply cr_left with (b := x).
    rewrite Heq ; apply le_refl.
    apply cr_trans with (U := U) ; auto.

    apply cr_left with (b := y).
    rewrite Heq ; apply le_refl.
    apply cr_trans with (U := W) ; auto.
  Qed.
  
  Lemma cov_inj_Covrel : forall U W, U ↪ W -> U ≤ W.
  Proof.
    intros.
    unfold le, Covrel_le, Covrel ; intros.
    unfold inclA in H.
    apply cr_refl. apply H. assumption.
  Qed.

  Ltac by_cov_inj :=
    try (apply cov_inj_Covrel) ;
    unfold inclA ;
    intro.

  Lemma covbij_coveq : forall U W : (list T), U == W -> U = W.
  Proof.
    intros.
    unfold equivlistA in H.
    split ; by_cov_inj ; intro ; apply H ; assumption.
  Qed.
  
  Lemma cr_right : forall a U W, a ◁ U -> U ↪ W -> a ◁ W.
  Proof.
    intros.
    apply cr_trans with (U := U).
    apply H.
    apply cov_inj_Covrel.
    apply H0.
  Qed.

  (** ** Binary join *)

  Instance CJoin : Join (list T) := (@app T).
  Ltac unfold_CJoin := unfold join, CJoin.

  Proposition CJoin_l : forall U V, U ≤ U ⊔ V.
  Proof.
    intros.
    by_cov_inj.
    unfold_CJoin.
    intros.
    rewrite InA_app_iff. left. assumption.
  Qed.

  Proposition CJoin_r : forall U V, V ≤ U ⊔ V.
  Proof.
    intros.
    by_cov_inj. unfold_CJoin. intros.
    rewrite InA_app_iff. right. assumption.
  Qed.

  Proposition CJoin_univ : forall U V W, U ≤ W -> V ≤ W ->
                                    U ⊔ V ≤ W.
  Proof.
    intros.
    unfold_CJoin. unfold_Covrel. intros.
    setoid_rewrite InA_app_iff in H1.
    destruct H1.
    apply H. assumption.
    apply H0. assumption.
  Qed.

  Add Morphism CJoin with signature (equiv_listT ==> equiv_listT ==> equiv_listT) as app_morphism.
  Proof.
    unfold equiv_listT, equivlistA. intros.
    unfold_CJoin. split ; intro ;
    setoid_rewrite InA_app_iff in H1 ;
    setoid_rewrite InA_app_iff.
    rewrite <- H, <- H0.
    assumption.
    rewrite H, H0.
    assumption.
  Qed.

  Lemma CJoin_comm : forall U V : list T, U ++ V == V ++ U.
  Proof.
    intros.
    unfold equivlistA. intros. split ; intros ; (
    setoid_rewrite InA_app_iff in H ;
    setoid_rewrite InA_app_iff ;
    destruct H ;
    [ right ; assumption |
      left ; assumption ]).
  Qed.

  (** We will get this fact for free from the
      distributive lattice structure we will define,
      but we need it before in the definition of the
      meet, so we prove it again here. *)

  Lemma CJoin_le_proper : Proper ((≤) ==> (≤) ==> (≤)) CJoin.
  Proof.
    unfold Proper, respectful.
    unfold_CJoin. intros.
    unfold_Covrel. intros.
    setoid_rewrite InA_app_iff in H1.
    destruct H1.
    - apply cr_right with (U := y).
      apply H. assumption.
      apply inclA_app_l.
    - apply cr_right with (U := y0).
      apply H0. assumption.
      apply inclA_app_r.
  Qed.

  (** Our temporary version of the finite joins: *)

  Definition Vl : list (list T) -> list T := @concat T.

  Lemma Vl_cons : forall u a, Vl (a :: u) = a ⊔ Vl u.
  Proof.
    intros. unfold_CJoin. unfold Vl.
    rewrite concat_cons.
    reflexivity.
  Qed.

  (** ** Binary meet *)
   
  Proposition cr_loc : forall a b U, a ◁ U -> b ⊓ a ◁ b ↓ U.
  Proof.
    intros a b U HR.
    induction HR as [a | a | a | a].

    - (* cr_bot *)
      rewrite H.
      meetsemilattice.
      simpl.
      apply cr_bot.
      reflexivity.
      
    - (* cr_refl *)
      apply cr_refl.
      unfold down ; simpl.
      apply map_in.
      unfold Proper, respectful. intros. rewrite H0. reflexivity.
      assumption.

    - (* cr_inf *)
      apply cr_inf with (b := b0) (i := i).
      apply le_trans with (y := a).
      apply meet_r. assumption.
      intros.
      rewrite <- meet_assoc.
      apply H1. assumption.

    - (* cr_left *)
      apply cr_left with (b := b ⊓ b0).
      apply meet_le_r ; assumption.
      apply IHHR.    
  Qed.

  Definition list_prod {A : Type} (f : T -> T -> A) (u v : list T) :=
    fold_left (fun accu x => accu ++ (map (f x) v)) u [].

  Lemma fold_left_concat : forall {A} (f : T -> T -> A) u v ac,
                             fold_left (fun accu x => accu ++ (map (f x) v)) u ac ≡ ac ++ (list_prod f u v).
  Proof.
    intros.
    generalize ac.
    induction u ; intros ; simpl.
    - rewrite app_nil_r. reflexivity.
    - unfold list_prod. simpl.
      rewrite IHu. rewrite IHu.
      rewrite app_assoc.
      reflexivity.
 Qed.
      
  Lemma list_prod_univ f : forall U V x, x ∈ (list_prod f U V) -> exists a b, a ∈ U /\ b ∈ V /\ x = f a b.
  Proof.
    intros.
    induction U ; simpl in H. inversion H.
    unfold list_prod in H. simpl in H.
    rewrite fold_left_concat in H.
    apply InA_app in H.
    destruct H.
    - apply in_map in H.
      destruct H as [y [H G]].
      exists a. exists y. split.
      + apply InA_cons_hd. reflexivity.
      + split ; assumption.
    - apply IHU in H.
      destruct H as (c & d & G & K & L).
      exists c. exists d. split.
      + apply InA_cons_tl. assumption.
      + split ; assumption.
  Qed.

  Lemma list_prod_inj f : Proper (Feq ==> Feq ==> Feq) f -> forall U V a b, a ∈ U -> b ∈ V -> (f a b) ∈ list_prod f U V.
  Proof.
    intros P U V a b H.
    generalize V. clear V.
    induction H ; intros V H' ;
    ( unfold list_prod ; simpl ;
      rewrite fold_left_concat ;
      setoid_rewrite InA_app_iff).
    - left.
      (* Quite tedious rewriting, I might be missing 
         an instance somewhere, but where? *)
      assert (f a b = f y b).
      apply P. assumption. reflexivity.
      set (Q := InA_Feq_compat).
      unfold Proper, respectful in Q.
      assert (equivlistA Feq (map (f y) V) (map (f y) V)) as K by reflexivity.
      specialize (Q (f a b) (f y b) H0 (map (f y) V) (map (f y) V) K).
      destruct Q.
      apply H2.
      apply map_in.
      apply P. reflexivity. assumption.
    - right.
      apply IHInA. assumption.
  Qed.
  
  Definition CMeet (U W : list T) : list T :=
    list_prod (⊓) U W.

  Instance CMeet_meet : Meet (list T) | 50 := CMeet.
  Ltac unfold_CMeet := unfold meet, CMeet_meet, CMeet.

  Proposition CMeet_l : forall U V : list T, U ⊓ V ≤ U.
  Proof.
    intros.
    unfold_CMeet.
    unfold_Covrel. intros.
    apply list_prod_univ in H.
    destruct H as (a & b & G & K & H).
    rewrite H.
    apply cr_left with (b := a).
    apply meet_l.
    apply cr_refl. assumption.
  Qed.

  Proposition CMeet_r : forall U V : list T, U ⊓ V ≤ V.
  Proof.
    intros.
    unfold_CMeet.
    unfold_Covrel. intros.
    apply list_prod_univ in H.
    destruct H as (a & b & G & K & H).
    rewrite H.
    apply cr_left with (b := b).
    apply meet_r.
    apply cr_refl. assumption.
  Qed.

  Lemma other_Covrel : forall U V : list T, U ≤ V <-> (forall x, x ◁ U -> x ◁ V).
  Proof.
    intros.
    split ; intros.
    - apply cr_trans with (U := U) ; assumption.
    - unfold_Covrel. intros.
      apply H. apply cr_refl. assumption.
  Qed.

  Lemma meet_elem_cov : forall U V x, x ∈ U -> map (x ⊓) V ↪ U ⊓ V.
  Proof.
    intros.
    induction H ; (
    unfold_CMeet ;
      unfold list_prod ; simpl ;
      rewrite fold_left_concat ;
      unfold inclA ; intros ;
      rewrite InA_app_iff).
    - left.
      assert (eqlistA Feq (map (x ⊓) V) (map (y ⊓) V)).
      clear H0.
      induction V. reflexivity.
      simpl. apply eqlistA_cons.
      rewrite H. reflexivity.
      apply IHV.
      rewrite <- H1.
      assumption.
    - right.
      apply IHInA. assumption.
  Qed.

  Lemma meet_covrel : forall x y U, y ◁ U -> x ⊓ y ◁ map (x ⊓) U.
  Proof.
    intros.
    induction H.
    - rewrite H. meetsemilattice.
      simpl.
      apply cr_bot. reflexivity.
    - apply cr_refl. apply map_in.
      apply meet_morphism_Proper. reflexivity.
      assumption.
    - apply cr_inf with (b := b) (i := i).
      apply le_trans with (y := a).
      apply meet_r. assumption.
      intros. rewrite <- meet_assoc.
      apply H1. assumption.
    - apply cr_left with (b := x ⊓ b).
      apply meet_le_r. assumption.
      assumption.
  Qed.

  Lemma CMeet_univ_internal : forall U V : list T, forall x y,
                                x ◁ U ->
                                y ◁ V ->
                                x ⊓ y ◁ U ⊓ V.
  Proof.
    intros.
    induction H.
    - rewrite H. meetsemilattice.
      apply cr_bot. reflexivity.
    - apply meet_elem_cov with (V := V) in H.
      apply cov_inj_Covrel in H.
      apply cr_trans with (U := map (a ⊓) V).
      apply meet_covrel. assumption.
      assumption.
    - apply cr_inf with (b := b) (i := i).
      apply le_trans with (y0 := a).
      apply meet_l. assumption.
      intros.
      rewrite <- meet_assoc.
      assert (y ⊓ x = x ⊓ y) by (apply meet_comm).
      rewrite H4.
      rewrite meet_assoc.
      apply H2. assumption.
    - apply cr_left with (b := b ⊓ y).
      apply meet_le_l. assumption.
      assumption.
  Qed.

  Proposition CMeet_univ : forall U V W : list T, W ≤ U -> W ≤ V -> W ≤ U ⊓ V.
  Proof.
    setoid_rewrite other_Covrel.
    intros.
    apply H0 in H1 as K.
    apply H in H1 as G.
    assert (x = x ⊓ x) by (rewrite meet_idem ; reflexivity).
    rewrite H2.
    apply CMeet_univ_internal ; assumption.
  Qed.

  (** ** Top and bottom *)

  Instance BotListT : Bottom (list T) := [].

  Lemma Bot_le : forall U, ⊥ ≤ U.
  Proof.
    intro.
    unfold_Covrel. intros.
    inversion H.
  Qed.

  Instance TopListT : Top (list T) := [ ⊤ ].
  Lemma Top_le : forall U : list T, U ≤ ⊤.
  Proof.
    intro.
    unfold_Covrel.
    intros.
    apply cr_left with (b := ⊤).
    apply top_le.
    apply cr_refl.
    apply InA_cons_hd.
    reflexivity.
  Qed.

  Instance MSL_for_FDistrLat : MeetSemiLattice Covrel :=
    MkMSL
      (list T)
      Covrel
      PO_for_FDistrLattice
      TopListT
      Top_le
      BotListT
      Bot_le
      CMeet
      CMeet_l
      CMeet_r
      CMeet_univ.
      

  (** ** Distributivity of binary meets over joins *)

  Lemma Cdistr_l : forall a b c, a ⊓ (b ⊔ c) ≤ (a ⊓ b) ⊔ (a ⊓ c).
  Proof.
    intros.
    (*assert (a ⊓ (b ⊔ c) = (b ⊔ c) ⊓ a) by (apply meet_comm).
    rewrite H. *)
    unfold meet, msl_meet, MSL_for_FDistrLat.
    unfold_CMeet.
    induction a ; unfold list_prod ; simpl.
    - simpl.
      apply Bot_le.
    - repeat (progress (rewrite fold_left_concat)).
      unfold join, CJoin.
      rewrite app_assoc.
      assert (forall w x y z : list T, (((w ++ x) ++ y) ++ z) = ((w ++ y) ++ (x ++ z))).
      + intros.
        apply covbij_coveq.
        assert ((w ++ x) ++ y == y ++ (w ++ x)) by (apply CJoin_comm).
        rewrite H.
        rewrite app_assoc. rewrite app_assoc.
        assert ((y ++ w) == (w ++ y)) by (apply CJoin_comm).
        rewrite H0.
        reflexivity.
      + rewrite H.
        apply CJoin_le_proper.
        * rewrite map_app.
          apply le_refl.
        * assumption.
  Qed.

  Instance FDistrLat : @DistrLattice (list T) Covrel :=
    MkDistrLattice
      (list T)
      Covrel
      MSL_for_FDistrLat
      CJoin
      CJoin_l
      CJoin_r
      CJoin_univ
      Cdistr_l.

  Definition LFeq := @Feq (list T) Covrel.
  Definition LFeq_setoid := Feq_equivalence PO_for_FDistrLattice.

  (** * Properties of the free distributive lattice *)
  
  (** ** Injection of generators *)

  Definition inj_gen (t : T) : (list T) := [t].

  Instance inj_gen_mslmorph : MSLMorphism Tmsl MSL_for_FDistrLat inj_gen.
  Proof.
    apply MkMSLMorphism ; unfold inj_gen.
    - apply MkPOMorphism.
      intros.
      unfold le, Covrel. intros.
      inversion H0.
      apply cr_left with (b := y).
      rewrite H2. assumption.
      apply cr_refl. apply InA_cons_hd. reflexivity.
      inversion H2.
    - intros.
      reflexivity.
    - split ; unfold_Covrel ; intros.
      + inversion H.
        rewrite H1.
        apply cr_bot. reflexivity.
        inversion H1.
      + inversion H.
    - reflexivity.
  Qed.
    
  Lemma V_inj_gen : forall u : list T, Vl (map inj_gen u) ≡ u.
  Proof.
    intro.
    induction u.
    - reflexivity.
    - simpl.
      rewrite IHu.
      reflexivity.
  Qed.
  
  Lemma inj_gen_le : forall t u, inj_gen t ≤ u <-> t ◁ u.
  Proof.
    intros.
    unfold inj_gen.
    unfold_Covrel.
    split ; intros.
    apply (H t).
    apply InA_cons_hd. reflexivity.
    inversion H0. subst.
    rewrite H2. assumption.
    inversion H2.
  Qed.

  Lemma inj_gen_meet : forall t u, inj_gen t ⊓ u = map (t ⊓) u.
  Proof.
    intros.
    reflexivity.
  Qed.

  (** ** Equalities generated by the axioms *)

  Proposition CovAx_meet_gen :
    forall (b:T), forall (i : Idx b), inj_gen b = (inj_gen b) ⊓ (CovAx b i).
  Proof.
    intros.
    rewrite inj_gen_meet.
    split.
    - rewrite inj_gen_le.
      apply cr_inf with (b := b) (i := i).
      apply le_refl.
      intros.
      apply cr_refl.
      apply map_in.
      + unfold Proper, respectful. intros.
        rewrite H0. reflexivity.
      + assumption.
    - rewrite <- inj_gen_meet.
      apply meet_l.
  Qed.

  Proposition CovAx_le_eq :
    forall (b:T), forall (i : Idx b), CovAx b i ≤ inj_gen b -> inj_gen b = CovAx b i.
  Proof.
    intros.
    split.
    - rewrite CovAx_meet_gen with (i := i).
      apply meet_r.
    - assumption.
  Qed.

  (** ** Universality *)
  
  (** Let us assume that we have a meet semilattice
     morphism to an arbitrary distributive lattice [R]. *)
  Context {R : Type}.
  Context {Rle : Le R}.
  Variable RDistrLat : @DistrLattice R Rle.

  Definition Rmsl := @dl_msl R Rle RDistrLat.
  Definition Rpo := @msl_preorder R Rle Rmsl.
  Variable f : T -> R.
  Variable mslmorph : MSLMorphism Tmsl Rmsl f.
  Existing Instance mslmorph.

  (** We assume that the morphism respects the axioms
      we have used to generate our free frame. *)
  Definition respects_axioms : Prop :=
    forall t : T, forall i : Idx t, f t ≤ Vf (map f (CovAx t i)).
  Variable resp_ax : respects_axioms.

  (** We define a function from our free frame to R. *)
  Definition fframe_ext (x : list T) : R :=
    Vf (map f x).

  (* We show that this function is a frame morphism. *)
  Existing Instance Covrel_le.

  (*
  Lemma f_covrel : forall a U, a ◁ U -> f a ≤ Vf (map f U).
  Proof.
    intros.
    induction H.
    - rewrite H.
      rewrite mslmorph_bot.
      apply @bot_le.
      exact mslmorph.
    - apply Vf_in_le.
      (* TODO *)

      rewrite <- H.
      assert (f (U n) = (f ∘ U) n) by reflexivity.
      rewrite H0 ; apply v_le.
    - unfold respects_axioms in resp_ax.
      specialize (resp_ax b i).
      set (K := (V (fun n => f (a ⊓ CovAx b i n)))).
      apply le_trans with (y := K).
      + assert (K = f a ⊓ V (f ∘ CovAx b i)).
        * rewrite cdistr.
          apply V_morphism ; intro.
          unfold compose.
          rewrite mslmorph_meet.
          reflexivity.
          apply mslmorph.
        * rewrite H2.
          apply le_trans with (y := f a ⊓ f b).
          assert (f a ≤ f b) by (apply (pomorph_le a b H)).
          assert (f a ⊓ f b = f a) by (apply order_meet ; assumption).
          rewrite H4.
          apply le_refl.
          apply meet_le.
          apply le_refl.
          assumption.
      + unfold K.
        apply v_univ.
        assumption.
    - apply le_trans with (y := f b).
      assert (f a ≤ f b) by (apply (pomorph_le a b H)).
      assumption. assumption.
  Qed.

  Instance fframe_mor : FMorphism FFrame RFrame fframe_ext.
  Proof.
    unfold fframe_ext.
    apply MkFMorphism.
    
    - apply MkMSLMorphism.
      + apply MkPOMorphism.
        intros.
        apply v_univ ; intro.
        unfold compose.
        unfold le, Covrel in H.
        specialize (H n).
        apply f_covrel ; assumption.
      + intros.
        unfold meet, msl_meet, FFrame. simpl.
        unfold CMeet, compose.
        assert (forall n, f (x (bijNN1 n) ⊓ y (bijNN2 n)) = f (x (bijNN1 n)) ⊓ f (y (bijNN2 n))).
        intro.
        apply (@mslmorph_meet T R Tle Rle Tmsl Rmsl f mslmorph).
        setoid_rewrite H.
        symmetry.
        apply V_meet.

      + unfold compose.
        unfold bottom, msl_bot, FFrame, Bot. simpl.
        assert (pointwise_relation nat Feq (fun _ => f ⊥) (fun _ => ⊥)).
        unfold pointwise_relation ; intro.
        apply mslmorph_bot. assumption.
        rewrite H.
        apply V_bot.

      + unfold compose.
        unfold top, msl_top, FFrame. simpl.
        rewrite V_top. reflexivity.
        exists O. unfold Top. apply mslmorph_top.
        apply mslmorph.

    - intro.
      unfold compose.
      rewrite <- V_pair.
      apply V_morphism ; intro.
      unfold V, FFrame, Vc, bijNN1, bijNN2.
      reflexivity.
  Qed.
  
  Definition fframe_mslmorph := fmorph_mslmorph FFrame RFrame fframe_ext.
  Proposition fframe_factoring : fframe_ext ∘ inj_gen = f.
  Proof.
    unfold equiv, ext_equiv, respectful.
    intros.
    unfold inj_gen, fframe_ext, compose.
    rewrite <- H.
    apply V_const.
  Qed.

  Arguments fframe_factoring : default implicits.

  (* Now the uniqueness part of the universality:
     if we have another such frame morphism,
     then it is equal to fframe_ext *)

  Variable other_fact : (list T) -> R.
  Variable other_morph : FMorphism FFrame RFrame other_fact.
  Existing Instance other_morph.
  Instance other_mslmorph : MSLMorphism MSL_for_FFrame Rmsl other_fact := fmorph_mslmorph FFrame RFrame other_fact.
  Instance other_morph_po : POMorphism other_fact.
  Proof.
    apply (mslmorph_pomorph MSL_for_FFrame Rmsl).
  Qed.    
    
  Variable other_commutes : other_fact ∘ inj_gen = f.

  Existing Instance Covrel_le.
  Instance coveq_R : Equiv (nat -> R) := @ext_equiv nat (≡) R (=).
  
  Proposition other_fact_equal : forall u, other_fact u = fframe_ext u.
  Proof.
    intro.
    assert (other_fact u = other_fact (V (fun n => inj_gen (u n)))).
    rewrite V_inj_gen ; reflexivity.
    rewrite H.
    rewrite morph_V.
    unfold fframe_ext, compose.
    apply V_morphism.
    intro.
    unfold equiv, ext_equiv, respectful in other_commutes.
    apply other_commutes ; reflexivity.
    assumption.
  Qed.
 *)
End Definition_Inductive_Locale.